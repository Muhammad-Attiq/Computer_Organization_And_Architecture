module KeypadScanner( 
    input [3:0] R,   
    input [2:0] C,   
    output [3:0] N,  
    output V         
); 
    assign N = (R == 4'b0001 && C == 3'b001) ? 4'b0001 :  
               (R == 4'b0001 && C == 3'b010) ? 4'b0010 :  
               (R == 4'b0001 && C == 3'b100) ? 4'b0011 :  
               (R == 4'b0010 && C == 3'b001) ? 4'b0100 :  
               (R == 4'b0010 && C == 3'b010) ? 4'b0101 :  
               (R == 4'b0010 && C == 3'b100) ? 4'b0110 :  
               (R == 4'b0100 && C == 3'b001) ? 4'b0111 :  
               (R == 4'b0100 && C == 3'b010) ? 4'b1000 :  
               (R == 4'b0100 && C == 3'b100) ? 4'b1001 :  
               (R == 4'b1000 && C == 3'b001) ? 4'b1010 :  
               (R == 4'b1000 && C == 3'b010) ? 4'b0000 :  
               (R == 4'b1000 && C == 3'b100) ? 4'b1011 :  
               4'b0000;  
 
    assign V = (R == 4'b0001 && (C == 3'b001 || C == 3'b010 || C == 3'b100)) || 
               (R == 4'b0010 && (C == 3'b001 || C == 3'b010 || C == 3'b100)) || 
               (R == 4'b0100 && (C == 3'b001 || C == 3'b010 || C == 3'b100)) || 
               (R == 4'b1000 && (C == 3'b001 || C == 3'b010 || C == 3'b100)); 
 
endmodule
